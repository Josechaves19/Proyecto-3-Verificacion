`include "uvm_macros.svh"
import uvm_pkg::*; 
`include "sequence_item.sv"
`include "sequence.sv"
`include "sequencer.sv"


module tb;

initial begin
    $display("HOlA"); 
    end
 endmodule

